// Copyright 2021 Thales DIS design services SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// Original Author: Guillaume Chauvon (guillaume.chauvon@thalesgroup.com)



package cvxif_instr_pkg;

  typedef enum logic [3:0] {
    LOAD_DENSE = 4'b0001,
    LOAD_SPARSE = 4'b0001,
    RESET_ACC = 4'b0001,
    STORE_ACC = 4'b0001,
  } opcode_t;


  typedef struct packed {
    logic accept;
    logic writeback;  // TODO depends on dualwrite
    logic [2:0] register_read;  // TODO Nr read ports
  } issue_resp_t;

  typedef struct packed {
    logic        accept;
    logic [31:0] instr;
  } compressed_resp_t;

  typedef struct packed {
    logic [31:0] instr;
    logic [31:0] mask;
    issue_resp_t resp;
    opcode_t     opcode;
  } copro_issue_resp_t;


  typedef struct packed {
    logic [15:0]      instr;
    logic [15:0]      mask;
    compressed_resp_t resp;
  } copro_compressed_resp_t;

  // 4 Possible RISCV instructions for Coprocessor
  parameter int unsigned NbInstr = 4;
  parameter copro_issue_resp_t CoproInstr[NbInstr] = '{
      '{
          // Custom LOAD DENSE
          instr:
          32'b00000_00_00000_00000_0_01_00000_0001011,  // custom0 opcode
          mask: 32'b11111_11_00000_00000_1_11_00000_1111111,
          resp : '{accept : 1'b1, writeback : 1'b0, register_read : {1'b0, 1'b1, 1'b1}},
          opcode : LOAD_DENSE
      },
      '{
          // Custom LOAD_SPARSE
          instr:
          32'b00000_00_00000_00000_0_10_00000_0001011,  // custom0 opcode
          mask: 32'b11111_11_00000_00000_1_11_00000_1111111,
          resp : '{accept : 1'b1, writeback : 1'b0, register_read : {1'b0, 1'b1, 1'b1}},
          opcode : LOAD_SPARSE
      },
      '{
          // Custom RESET_ACC
          instr:
          32'b00000_01_00000_00000_0_00_00000_0001011,  // custom0 opcode
          mask: 32'b11111_11_00000_00000_1_11_00000_1111111,
          resp : '{accept : 1'b1, writeback : 1'b0, register_read : {1'b0, 1'b0, 1'b0}},
          opcode : RESET_ACC
      },
      '{
          // Custom STORE_ACC
          instr:
          32'b00000_10_00000_00000_0_11_00000_0001011,  // custom0 opcode
          mask: 32'b11111_11_00000_00000_1_11_00000_1111111,
          resp : '{accept : 1'b1, writeback : 1'b1, register_read : {1'b0, 1'b0, 1'b1}},
          opcode : STORE_ACC
      }
  };

endpackage
